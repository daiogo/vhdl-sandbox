library verilog;
use verilog.vl_types.all;
entity hamming_weight_calculator_vlg_vec_tst is
end hamming_weight_calculator_vlg_vec_tst;
