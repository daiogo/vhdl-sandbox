library verilog;
use verilog.vl_types.all;
entity signed_adder_vlg_vec_tst is
end signed_adder_vlg_vec_tst;
