library verilog;
use verilog.vl_types.all;
entity arbiter_vlg_vec_tst is
end arbiter_vlg_vec_tst;
