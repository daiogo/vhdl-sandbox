library verilog;
use verilog.vl_types.all;
entity code_converter_vlg_vec_tst is
end code_converter_vlg_vec_tst;
