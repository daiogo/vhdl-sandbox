library verilog;
use verilog.vl_types.all;
entity reference_setter_vlg_vec_tst is
end reference_setter_vlg_vec_tst;
