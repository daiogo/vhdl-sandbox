library verilog;
use verilog.vl_types.all;
entity multiple_detector_vlg_vec_tst is
end multiple_detector_vlg_vec_tst;
