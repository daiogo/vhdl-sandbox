library verilog;
use verilog.vl_types.all;
entity password_detector_vlg_vec_tst is
end password_detector_vlg_vec_tst;
