library verilog;
use verilog.vl_types.all;
entity decoder_3to2_vlg_vec_tst is
end decoder_3to2_vlg_vec_tst;
