library verilog;
use verilog.vl_types.all;
entity random_onehot_generator_vlg_vec_tst is
end random_onehot_generator_vlg_vec_tst;
