library verilog;
use verilog.vl_types.all;
entity pseudorandom_generator_vlg_vec_tst is
end pseudorandom_generator_vlg_vec_tst;
