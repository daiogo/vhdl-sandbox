library verilog;
use verilog.vl_types.all;
entity tflipflop_vlg_vec_tst is
end tflipflop_vlg_vec_tst;
