library verilog;
use verilog.vl_types.all;
entity synchronous_counter_vlg_vec_tst is
end synchronous_counter_vlg_vec_tst;
